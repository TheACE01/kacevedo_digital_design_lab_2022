module vga_controller(
	input logic clk,
	input logic rst,
	input logic VGA_CLK,
	input logic [9:0] h_counter, v_counter,
	output logic VGA_HS,
	output logic VGA_VS,
	output logic VGA_BLANK_N,
	output logic VGA_SYNC_N,
	output logic video_on);				
    
    // 800 pixels per line (including front/back porch)
    // 525 lines per frame (including front/back porch)
    parameter [9:0] H_TOTAL = 10'd800;
    parameter [9:0] V_TOTAL = 10'd525;
    
    logic VGA_HS_in, VGA_VS_in, VGA_BLANK_N_in;
    assign VGA_SYNC_N = 1'b0;
	 
	 // Define the video on signal
	 assign video_on = VGA_BLANK_N;
    
    // VGA control signals. 
    // VGA_CLK is generated by PLL
    always_ff @ (posedge VGA_CLK or negedge rst) begin
        if (!rst) begin
            VGA_HS <= 1'b0;
            VGA_VS <= 1'b0;
            VGA_BLANK_N <= 1'b0;
        end
        else begin
            VGA_HS <= VGA_HS_in;
            VGA_VS <= VGA_VS_in;
            VGA_BLANK_N <= VGA_BLANK_N_in;
        end
    end
	 
    
    always_comb begin
        // Horizontal sync pulse is 96 pixels long at pixels 656-752
        VGA_HS_in = 1'b1;
        if(h_counter >= 10'd656 && h_counter < 10'd752)
            VGA_HS_in = 1'b0;
				
        // Vertical sync pulse is 2 lines (800 pixels each) long at line 490-491
        VGA_VS_in = 1'b1;
        if(v_counter >= 10'd490 && v_counter < 10'd492)
            VGA_VS_in = 1'b0;
				
        // Display pixels (inhibit blanking) between horizontal 0-639 and vertical 0-479 (640x480)
        VGA_BLANK_N_in = 1'b0;
        if(h_counter < 10'd640 && v_counter < 10'd480)
            VGA_BLANK_N_in = 1'b1;
    end
endmodule
