module deco_binario_bcd (A3, A2, A1, A0, S4, S3, S2, S1, S0);

  input logic A3, A2, A1, A0;
  output logic S4, S3, S2, S1, S0;
  
  
endmodule
